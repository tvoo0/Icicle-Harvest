`timescale 1ns / 1ps

module hex7seg(
     input [3:0] n,
     input negative,
     output [6:0] seg
    );
    
    assign seg[0] = negative | (~n[3]&~n[2]&~n[1]&n[0])|(~n[3]&n[2]&~n[1]*~n[0])|(n[3]&~n[2]&n[1]&n[0])|(n[3]&n[2]&~n[1]&n[0]);
    assign seg[1] = negative | (~n[3]&n[2]&~n[1]&n[0])|(~n[3]&n[2]&n[1]&~n[0])|(n[3]&~n[2]&n[1]&n[0])|(n[3]&n[2]&~n[1]&~n[0])|(n[3]&n[2]&n[1]&~n[0])|(n[3]&n[2]&n[1]&n[0]);
    assign seg[2] = negative | (~n[3]&~n[2]&n[1]&~n[0])|(n[3]&n[2]&~n[1]&~n[0])|(n[3]&n[2]&n[1]&~n[0])|(n[3]&n[2]&n[1]&n[0]);
    assign seg[3] = negative | (~n[3]&~n[2]&~n[1]&n[0])|(~n[3]&n[2]&~n[1]&~n[0])|(~n[3]&n[2]&n[1]&n[0])|(n[3]&~n[2]&~n[1]&n[0])|(n[3]&~n[2]&n[1]&~n[0])|(n[3]&n[2]&n[1]&n[0]);
    assign seg[4] = negative | (~n[3]&~n[2]&~n[1]&n[0])|(~n[3]&~n[2]&n[1]&n[0])|(~n[3]&n[2]&~n[1]&~n[0])|(~n[3]&n[2]&~n[1]&n[0])|(~n[3]&n[2]&n[1]&n[0])|(n[3]&~n[2]&~n[1]&n[0]);
    assign seg[5] = negative | (~n[3]&~n[2]&~n[1]&n[0])|(~n[3]&~n[2]&n[1]&~n[0])|(~n[3]&~n[2]&n[1]&n[0])|(~n[3]&n[2]&n[1]&n[0])|(n[3]&n[2]&~n[1]&n[0]);
    assign seg[6] = ~negative & (~n[3]&~n[2]&~n[1]&~n[0])|(~n[3]&~n[2]&~n[1]&n[0])|(~n[3]&n[2]&n[1]&n[0])|(n[3]&n[2]&~n[1]&~n[0]);
    
endmodule